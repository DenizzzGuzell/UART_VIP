package uart_agent_pkg_tx;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "../../../utils/config_macro.svh"
	
	`include "uart_seq_item_tx.svh"
	`include "uart_sequencer_tx.svh"
	`include "uart_agent_config_tx.svh"
	`include "uart_driver_tx.svh"
	`include "uart_monitor_tx.svh"
	`include "uart_agent_tx.svh"
	
endpackage: uart_agent_pkg_tx