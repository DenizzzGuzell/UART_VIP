package uart_agent_pkg_rx;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "../../../utils/config_macro.svh"

	`include "uart_seq_item_rx.svh"
	`include "uart_sequencer_rx.svh"
	`include "uart_agent_config_rx.svh"
	`include "uart_driver_rx.svh"
	`include "uart_monitor_rx.svh"
	`include "uart_agent_rx.svh"

endpackage: uart_agent_pkg_rx
